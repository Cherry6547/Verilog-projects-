module EighttoThreeEncoder_tb;
    reg [7:0]a;
    wire [0:2]y;
    EighttoThreeEncoder uut(
        .a(a),
        .y(y)
    );
    initial begin
        $dumpfile("EighttoThreeEncoder.vcd");
        $dumpvars(0,EighttoThreeEncoder_tb);
        a = 8'b00000001;
        #10 a = 8'b00000010;
        #10 a = 8'b00000100;
        #10 a = 8'b00001000;
        #10 a = 8'b00010000;
        #10 a = 8'b00100000;
        #10 a = 8'b01000000;
        #10 a = 8'b10000000;
        #10 $finish;
    end
endmodule