module BcdtoXs3(
    input [3:0]a,
    output [3:0]y
);
assign y = a + 3;
endmodule